module main();
    initial $display("Hello, World!");
endmodule
